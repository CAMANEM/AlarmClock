// cpu_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module cpu_tb (
	);

	wire        cpu_inst_clk_bfm_clk_clk;       // cpu_inst_clk_bfm:clk -> [cpu_inst:clk_clk, cpu_inst_reset_bfm:clk]
	wire  [1:0] cpu_inst_leds_export;           // cpu_inst:leds_export -> cpu_inst_leds_bfm:sig_export
	wire        cpu_inst_reset_bfm_reset_reset; // cpu_inst_reset_bfm:reset -> cpu_inst:reset_reset_n

	cpu cpu_inst (
		.clk_clk       (cpu_inst_clk_bfm_clk_clk),       //   clk.clk
		.leds_export   (cpu_inst_leds_export),           //  leds.export
		.reset_reset_n (cpu_inst_reset_bfm_reset_reset)  // reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) cpu_inst_clk_bfm (
		.clk (cpu_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm cpu_inst_leds_bfm (
		.sig_export (cpu_inst_leds_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) cpu_inst_reset_bfm (
		.reset (cpu_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (cpu_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
